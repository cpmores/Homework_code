/******************************************************************************
 ** Logisim-evolution goes FPGA automatic generated Verilog code             **
 ** https://github.com/logisim-evolution/                                    **
 **                                                                          **
 ** Component : logisimTopLevelShell                                         **
 **                                                                          **
 *****************************************************************************/

module logisimTopLevelShell(  );

   /*******************************************************************************
   ** The wires are defined here                                                 **
   *******************************************************************************/
   wire s_D;
   wire s_Q;
   wire s_Qbar;
   wire s_clk;
   wire s_mid_Q;

   /*******************************************************************************
   ** The module functionality is described here                                 **
   *******************************************************************************/

   /*******************************************************************************
   ** All signal adaptations are performed here                                  **
   *******************************************************************************/
   assign s_D   = 1'b0;
   assign s_clk = 1'b0;

   /*******************************************************************************
   ** The toplevel component is connected here                                   **
   *******************************************************************************/
   ms_sr_flip_flop   CIRCUIT_0 (.D(s_D),
                                .Q(s_Q),
                                .Qbar(s_Qbar),
                                .clk(s_clk),
                                .mid_Q(s_mid_Q));
endmodule
